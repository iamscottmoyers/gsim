-- Comment for a test vhdl file :)
entity a is
        port (l : in std_logic;
              art : out moosetype);
end

architecture tootle of a is
        begin
        end architecture tooTle;
entity b is
begin end
entity c is
begin end entity c
entity d is
begin end d
entity e is
begin end entity
